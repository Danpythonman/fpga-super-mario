module VgaCoin
(
	input [31:0] x,
	input [31:0] y,
	input byte background [11:0][16:0],
	input [3:0] background_red,
	input [3:0] background_green,
	input [3:0] background_blue,
	output reg [3:0] red,
	output reg [3:0] green,
	output reg [3:0] blue
);

	localparam NULL = 0;
	localparam COLOR1 = 1;
	localparam COLOR2 = 2;
	localparam COLOR3 = 3;
	localparam COLOR4 = 4;
	localparam COLOR5 = 5;
	localparam COLOR6 = 6;
	localparam COLOR7 = 7;
	localparam COLOR8 = 8;
	localparam COLOR9 = 9;
	localparam COLOR10 = 10;
	localparam COLOR11 = 11;
	localparam COLOR12 = 12;
	localparam COLOR13 = 13;
	localparam COLOR14 = 14;
	localparam COLOR15 = 15;
	localparam COLOR16 = 16;

	reg [5:0] pattern [38:0][38:0] = '{
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR4,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR4,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR4,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR4,
			COLOR2,
			COLOR2,
			COLOR2,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR2,
			COLOR2,
			COLOR2,
			COLOR2,
			COLOR2,
			COLOR2,
			COLOR2,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR2,
			COLOR5,
			COLOR6,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR3,
			COLOR3,
			COLOR4,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR3,
			COLOR3,
			COLOR3,
			NULL,
			NULL,
			COLOR6,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR3,
			COLOR3,
			COLOR4,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR6,
			COLOR6,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR3,
			COLOR3,
			COLOR2,
			NULL,
			NULL
		},
		'{
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR4,
			NULL,
			NULL,
			COLOR7,
			COLOR7,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR7,
			COLOR7,
			COLOR3,
			COLOR3,
			COLOR2,
			NULL,
			NULL
		},
		'{
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR4,
			NULL,
			COLOR9,
			COLOR7,
			COLOR7,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR7,
			COLOR7,
			COLOR3,
			COLOR3,
			COLOR4,
			NULL,
			NULL
		},
		'{
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR7,
			COLOR7,
			COLOR8,
			COLOR8,
			COLOR11,
			NULL,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			COLOR9,
			NULL,
			COLOR6,
			COLOR7,
			COLOR7,
			COLOR10,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3
		},
		'{
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR7,
			COLOR7,
			COLOR8,
			COLOR8,
			COLOR9,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR9,
			COLOR7,
			COLOR7,
			COLOR12,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3
		},
		'{
			COLOR2,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR13,
			COLOR7,
			COLOR7,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR11,
			COLOR6,
			COLOR6,
			COLOR6,
			COLOR6,
			COLOR2,
			COLOR14,
			COLOR15,
			COLOR7,
			COLOR7,
			COLOR12,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3
		},
		'{
			COLOR3,
			COLOR3,
			NULL,
			NULL,
			COLOR6,
			COLOR7,
			COLOR7,
			NULL,
			NULL,
			COLOR11,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR7,
			COLOR7,
			COLOR12,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3
		},
		'{
			COLOR3,
			COLOR3,
			COLOR2,
			NULL,
			COLOR6,
			COLOR7,
			COLOR7,
			NULL,
			NULL,
			COLOR11,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR7,
			COLOR7,
			COLOR12,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3
		},
		'{
			COLOR3,
			COLOR3,
			COLOR2,
			NULL,
			COLOR6,
			COLOR7,
			COLOR7,
			NULL,
			NULL,
			COLOR6,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR7,
			COLOR7,
			COLOR12,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3
		},
		'{
			COLOR3,
			COLOR3,
			NULL,
			NULL,
			COLOR6,
			COLOR7,
			COLOR7,
			NULL,
			NULL,
			COLOR6,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR7,
			COLOR7,
			COLOR12,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3
		},
		'{
			COLOR3,
			COLOR3,
			COLOR4,
			COLOR14,
			COLOR15,
			COLOR7,
			COLOR7,
			COLOR11,
			COLOR11,
			COLOR13,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR10,
			COLOR10,
			COLOR13,
			COLOR7,
			COLOR7,
			COLOR12,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3
		},
		'{
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR7,
			COLOR7,
			COLOR8,
			COLOR8,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR7,
			COLOR7,
			COLOR12,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3
		},
		'{
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR7,
			COLOR7,
			COLOR8,
			COLOR8,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR7,
			COLOR7,
			COLOR10,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3
		},
		'{
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR12,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR7,
			COLOR7,
			COLOR13,
			COLOR12,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR4,
			NULL,
			NULL
		},
		'{
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR12,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR7,
			COLOR7,
			COLOR13,
			COLOR10,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR2,
			NULL,
			NULL
		},
		'{
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR13,
			COLOR13,
			COLOR13,
			COLOR13,
			COLOR7,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR8,
			COLOR13,
			COLOR13,
			COLOR12,
			COLOR10,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR4,
			NULL,
			NULL
		},
		'{
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR13,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR12,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR2,
			NULL,
			NULL
		},
		'{
			NULL,
			COLOR2,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR13,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR7,
			COLOR12,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR2,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR12,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR10,
			COLOR12,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR10,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR2,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR3,
			COLOR16,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR16,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR4,
			COLOR2,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			COLOR3,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		},
		'{
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL,
			NULL
		}
	};

	always @(x, y) begin
		if (pattern[x][y] == NULL) begin
			red   <= background_red;
			green <= background_green;
			blue  <= background_blue;
		end else if (pattern[x][y] == COLOR1) begin
			red   <= 4'd13;
			green <= 4'd13;
			blue  <= 4'd13;
		end else if (pattern[x][y] == COLOR2) begin
			red   <= 4'd9;
			green <= 4'd9;
			blue  <= 4'd9;
		end else if (pattern[x][y] == COLOR3) begin
			red   <= 4'd2;
			green <= 4'd2;
			blue  <= 4'd2;
		end else if (pattern[x][y] == COLOR4) begin
			red   <= 4'd6;
			green <= 4'd6;
			blue  <= 4'd6;
		end else if (pattern[x][y] == COLOR5) begin
			red   <= 4'd9;
			green <= 4'd9;
			blue  <= 4'd13;
		end else if (pattern[x][y] == COLOR6) begin
			red   <= 4'd13;
			green <= 4'd9;
			blue  <= 4'd6;
		end else if (pattern[x][y] == COLOR7) begin
			red   <= 4'd13;
			green <= 4'd9;
			blue  <= 4'd2;
		end else if (pattern[x][y] == COLOR8) begin
			red   <= 4'd13;
			green <= 4'd13;
			blue  <= 4'd2;
		end else if (pattern[x][y] == COLOR9) begin
			red   <= 4'd13;
			green <= 4'd13;
			blue  <= 4'd9;
		end else if (pattern[x][y] == COLOR10) begin
			red   <= 4'd6;
			green <= 4'd6;
			blue  <= 4'd2;
		end else if (pattern[x][y] == COLOR11) begin
			red   <= 4'd13;
			green <= 4'd13;
			blue  <= 4'd6;
		end else if (pattern[x][y] == COLOR12) begin
			red   <= 4'd9;
			green <= 4'd6;
			blue  <= 4'd2;
		end else if (pattern[x][y] == COLOR13) begin
			red   <= 4'd9;
			green <= 4'd9;
			blue  <= 4'd2;
		end else if (pattern[x][y] == COLOR14) begin
			red   <= 4'd6;
			green <= 4'd6;
			blue  <= 4'd9;
		end else if (pattern[x][y] == COLOR15) begin
			red   <= 4'd9;
			green <= 4'd9;
			blue  <= 4'd6;
		end else if (pattern[x][y] == COLOR16) begin
			red   <= 4'd6;
			green <= 4'd2;
			blue  <= 4'd2;
		end	end

endmodule
